library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

ENTITY counter IS
	PORT (
		CLK : in  STD_LOGIC;
		RST : in  STD_LOGIC;
		O   : out STD_LOGIC_VECTOR( 7 DOWNTO 0)
	);
END counter;

ARCHITECTURE Behavioral OF counter IS
	SIGNAL COUNTER : UNSIGNED(7 DOWNTO 0);
BEGIN

	PROCESS(RST, CLK)
	BEGIN
		IF RST = '1' THEN
			COUNTER <= TO_UNSIGNED( 0, 8 );
		ELSIF CLK = '1' AND CLK'EVENT THEN
			COUNTER <= TO_UNSIGNED( 0, 8 );
		END IF;
	END PROCESS;

	O <= STD_LOGIC_VECTOR( COUNTER );

END Behavioral;